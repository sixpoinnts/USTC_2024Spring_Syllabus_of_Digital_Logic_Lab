module Shifter1(
    input                   [31 : 0]        src0,
    input                   [ 4 : 0]        src1,
    output     reg          [31 : 0]        res1,       //逻辑右移
    output     reg          [31 : 0]        res2        //算术右移
);
// Write your code here
always @(*) begin
    case (src1)
        5'd0:begin
            res1=src0;
            res2=src0;
        end 
        5'd1:begin
            res1={1'b0,src0[31:1]};
            res2={{1{src0[31]}},src0[31:1]};
        end 
        5'd2:begin
            res1={2'b0,src0[31:2]};
            res2={{2{src0[31]}},src0[31:2]};
        end 
        5'd3:begin
            res1={3'b0,src0[31:3]};
            res2={{3{src0[31]}},src0[31:3]};
        end 
        5'd4:begin
            res1={4'b0,src0[31:4]};
            res2={{4{src0[31]}},src0[31:4]};
        end 
        5'd5:begin
            res1={5'b0,src0[31:5]};
            res2={{5{src0[31]}},src0[31:5]};
        end 
        5'd6:begin
            res1={6'b0,src0[31:6]};
            res2={{6{src0[31]}},src0[31:6]};
        end 
        5'd7:begin
            res1={7'b0,src0[31:7]};
            res2={{7{src0[31]}},src0[31:7]};
        end 
        5'd8:begin
            res1={8'b0,src0[31:8]};
            res2={{8{src0[31]}},src0[31:8]};
        end 
        5'd9:begin
            res1={9'b0,src0[31:9]};
            res2={{9{src0[31]}},src0[31:9]};
        end 
        5'd10:begin
            res1={10'b0,src0[31:10]};
            res2={{10{src0[31]}},src0[31:10]};
        end 
        5'd11:begin
            res1={11'b0,src0[31:11]};
            res2={{11{src0[31]}},src0[31:11]};
        end 
        5'd12:begin
            res1={12'b0,src0[31:12]};
            res2={{12{src0[31]}},src0[31:12]};
        end 
        5'd13:begin
            res1={13'b0,src0[31:13]};
            res2={{13{src0[31]}},src0[31:13]};
        end 
        5'd14:begin
            res1={14'b0,src0[31:14]};
            res2={{14{src0[31]}},src0[31:14]};
        end 
        5'd15:begin
            res1={15'b0,src0[31:15]};
            res2={{15{src0[31]}},src0[31:15]};
        end 
        5'd16:begin
            res1={16'b0,src0[31:16]};
            res2={{16{src0[31]}},src0[31:16]};
        end 
        5'd17:begin
            res1={17'b0,src0[31:17]};
            res2={{17{src0[31]}},src0[31:17]};
        end 
        5'd18:begin
            res1={18'b0,src0[31:18]};
            res2={{18{src0[31]}},src0[31:18]};
        end 
        5'd19:begin
            res1={19'b0,src0[31:19]};
            res2={{19{src0[31]}},src0[31:19]};
        end 
        5'd20:begin
            res1={20'b0,src0[31:20]};
            res2={{20{src0[31]}},src0[31:20]};
        end 
        5'd21:begin
            res1={21'b0,src0[31:21]};
            res2={{21{src0[31]}},src0[31:21]};
        end 
        5'd22:begin
            res1={22'b0,src0[31:22]};
            res2={{22{src0[31]}},src0[31:22]};
        end 
        5'd23:begin
            res1={23'b0,src0[31:23]};
            res2={{23{src0[31]}},src0[31:23]};
        end 
        5'd24:begin
            res1={24'b0,src0[31:24]};
            res2={{24{src0[31]}},src0[31:24]};
        end 
        5'd25:begin
            res1={25'b0,src0[31:25]};
            res2={{25{src0[31]}},src0[31:25]};
        end 
        5'd26:begin
            res1={26'b0,src0[31:26]};
            res2={{26{src0[31]}},src0[31:26]};
        end 
        5'd27:begin
            res1={27'b0,src0[31:27]};
            res2={{27{src0[31]}},src0[31:27]};
        end 
        5'd28:begin
            res1={28'b0,src0[31:28]};
            res2={{28{src0[31]}},src0[31:28]};
        end 
        5'd29:begin
            res1={29'b0,src0[31:29]};
            res2={{29{src0[31]}},src0[31:29]};
        end 
        5'd30:begin
            res1={30'b0,src0[31:30]};
            res2={{30{src0[31]}},src0[31:30]};
        end 
        5'd31:begin
            res1={31'b0,src0[31]};
            res2={{31{src0[31]}},src0[31]};
        end 
    endcase
end
// End of your code
endmodule
