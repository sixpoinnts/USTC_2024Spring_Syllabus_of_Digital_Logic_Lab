module Uart_test (
    input                   [ 0 : 0]            uart_din,
    output                  [ 0 : 0]            uart_dout
);
assign uart_dout = uart_din;
endmodule
